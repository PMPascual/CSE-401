`timescale 1ns / 1ps

module Mem(
   output reg [31:0] data,      
   input wire [31:0] addr   
   );

   reg [31:0] MEM[0:127];
   integer i;

   // initial begin
   // MEM[0] <= 'bA00000AA;
   // MEM[1] <= 'b10000011;
   // MEM[2] <= 'b20000022;
   // MEM[3] <= 'b30000033;
   // MEM[4] <= 'b40000044;
   // MEM[5] <= 'b50000055;
   // MEM[6] <= 'b60000066;
   // MEM[7] <= 'b70000077;
   // MEM[8] <= 'b80000088;
   // MEM[9] <= 'b90000099;
   // end

   initial begin
   MEM[0] <= 'b10001100000000010000000000000001;
   MEM[1] <= 'b10001100000000010000000000000010;
   MEM[2] <= 'b10001100000000010000000000000011;
   MEM[3] <= 'b10000000000000000000000000000000;
   MEM[4] <= 'b10000000000000000000000000000000;
   MEM[5] <= 'b00000000001000100000100000100000;
   MEM[6] <= 'b10000000000000000000000000000000;
   MEM[7] <= 'b10000000000000000000000000000000;
   MEM[8] <= 'b10000000000000000000000000000000;
   MEM[9] <= 'b00000000001000110000100000100000;
   MEM[10] <= 'b10000000000000000000000000000000;
   MEM[11] <= 'b10000000000000000000000000000000;
   MEM[12] <= 'b10000000000000000000000000000000;
   MEM[13] <= 'b00000000001000010000100000100000;
   MEM[14] <= 'b10000000000000000000000000000000;
   MEM[15] <= 'b10000000000000000000000000000000;
   MEM[16] <= 'b10000000000000000000000000000000;
   MEM[17] <= 'b10000000000000000000000000000000;
   MEM[18] <= 'b00000000001000000000100000100000;
   MEM[19] <= 'b10000000000000000000000000000000;
   MEM[20] <= 'b10000000000000000000000000000000;
   MEM[21] <= 'b10000000000000000000000000000000;
   MEM[22] <= 'b10000000000000000000000000000000;
   MEM[23] <= 'b10000000000000000000000000000000;
   end
   
   // initial
   // $readmemb("/home/csusb.edu/005705423/Documents/risc.txt",MEM);
   // begin


   always @(addr) begin
		data <= MEM[addr];
   end
endmodule
